* D:\Project\project2.sch

* Schematics Version 9.2
* Wed Aug 31 15:22:04 2022



** Analysis setup **
.tran 10u 0.8 0.6 100u
.OP 
.LIB "D:\Project\project2.lib"


* From [PSPICE NETLIST] section of d:\orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "project2.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
